`timescale 1ns/1ps
`default_nettype none

module ovo7670_top
    #(

    ) (
        input wire clk_i, reset_i
    );

endmodule
