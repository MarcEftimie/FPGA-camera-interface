`timescale 1ns/1ps
`default_nettype none

module ovo7670_interface
    #(
    ) (
        input wire pclk_cmos_i, reset_i,
        input wire vsync_cmos_i,
        input wire href_cmos_i,
        output wire hsync_o
    );



endmodule
